* Spice output from KLayout SiEPIC-Tools v0.3.73, 2021-03-27 20:18:31.

.subckt test_mzi ebeam_gc_te1550_laser1 ebeam_gc_te1550_detector2
.param MC_uniformity_width=0 
.param MC_uniformity_thickness=0 
.param MC_resolution_x=100 
.param MC_resolution_y=100 
.param MC_grid=10e-6 
.param MC_non_uniform=99 
 ebeam_y_1550_0  N$0 N$1 N$2 ebeam_y_1550 library="Design kits/ebeam"  lay_x=-41.0E-6 lay_y=16.19E-6 sch_x=-3.591240876E0 sch_y=1.41810219E0 
 ebeam_gc_te1550_1  ebeam_gc_te1550_laser1 N$0 ebeam_gc_te1550 library="Design kits/ebeam"  lay_x=-64.9E-6 lay_y=16.19E-6 sch_x=-5.684671533E0 sch_y=1.41810219E0 
 ebeam_gc_te1550_2  ebeam_gc_te1550_detector2 N$3 ebeam_gc_te1550 library="Design kits/ebeam"  lay_x=-64.9E-6 lay_y=143.19E-6 sch_x=-5.684671533E0 sch_y=12.542189781E0 
 ebeam_y_1550_3  N$3 N$5 N$4 ebeam_y_1550 library="Design kits/ebeam"  lay_x=-41.0E-6 lay_y=143.19E-6 sch_x=-3.591240876E0 sch_y=12.542189781E0 
 ebeam_wg_integral_1550_4  N$1 N$4 ebeam_wg_integral_1550 library="Design kits/EBeam" wg_length=159.537u wg_width=0.500u points="[[-33.6,18.94],[-13.03,18.94],[-13.03,140.44],[-33.6,140.44]]" radius=5.0 lay_x=-22.94E-6 lay_y=79.69E-6 sch_x=-2.009343066E0 sch_y=6.980145985E0 
 ebeam_wg_integral_1550_5  N$5 N$2 ebeam_wg_integral_1550 library="Design kits/EBeam" wg_length=197.937u wg_width=0.500u points="[[-33.6,145.94],[0.67,145.94],[0.67,13.44],[-33.6,13.44]]" radius=5.0 lay_x=-16.09E-6 lay_y=79.69E-6 sch_x=-1.409343066E0 sch_y=6.980145985E0 
.ends test_mzi

test_mzi   ebeam_gc_te1550_laser1 ebeam_gc_te1550_detector2 test_mzi sch_x=-1 sch_y=-1 

* Spice output from KLayout SiEPIC-Tools v0.3.73, 2021-03-27 20:18:31.

* Optical Network Analyzer:
.ona input_unit=wavelength input_parameter=start_and_stop
  + minimum_loss=80
  + analysis_type=scattering_data
  + multithreading=user_defined number_of_threads=1
  + orthogonal_identifier=1
  + start=1500.000e-9
  + stop=1600.000e-9
  + number_of_points=2000
  + input(1)=test_mzi,ebeam_gc_te1550_detector2
  + output=test_mzi,ebeam_gc_te1550_laser1
.INCLUDE "C:\Users\jai\AppData\Local\Temp\tmpkij35j69\test_mzi.spi"

